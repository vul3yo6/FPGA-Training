`timescale 10ns / 1ps
module HA(s, c, x, y);
input x, y;
output s, c;

/*
    write your code here
*/

endmodule
