`timescale 10ns / 1ps
`include "FA.v"
module RCA(s, cout, x, y, c0);
input  [3:0] x, y;
output [3:0] s;
input  c0;
output cout;
wire c1, c2, c3;

/*
    write your code here
*/

endmodule
