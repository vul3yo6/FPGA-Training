`timescale 10ns / 1ps
`include "HA.v"
module FA(s, c_out, x, y, c_in);
input x, y, c_in;
output s, c_out;
wire s1, c1, c2;

/*
    write your code here
*/
  
endmodule

