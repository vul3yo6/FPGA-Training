`include "FA.v"
module AS(sel, A, B, S, O);
input [3:0] A, B;
input sel;
output [3:0] S;
output O;

/*
    write your code here
*/

endmodule


